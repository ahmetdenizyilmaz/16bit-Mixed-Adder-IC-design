*** SPICE deck for cell Or2Gate{sch} from library 16BitAdder
*** Created on Pzt Oca 07, 2019 17:16:27
*** Last revised on Paz Oca 13, 2019 20:38:34
*** Written on Paz Oca 13, 2019 20:54:11 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT _16BitAdder__Inverter FROM CELL Inverter{sch}
.SUBCKT _16BitAdder__Inverter Out Inp
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 Out Inp gnd gnd NMOS L=0.6U W=1.8U
Mpmos@1 vdd Inp Out vdd PMOS L=0.6U W=3.6U
.ENDS _16BitAdder__Inverter

*** SUBCIRCUIT _16BitAdder__Nor2Gate FROM CELL Nor2Gate{sch}
.SUBCKT _16BitAdder__Nor2Gate Out Inp0 Inp1
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Out Inp0 gnd gnd NMOS L=0.6U W=1.8U
Mnmos@1 Out Inp1 gnd gnd NMOS L=0.6U W=1.8U
Mpmos@0 net@11 Inp1 Out vdd PMOS L=0.6U W=3.6U
Mpmos@1 vdd Inp0 net@11 vdd PMOS L=0.6U W=3.6U
.ENDS _16BitAdder__Nor2Gate

.global gnd vdd

*** TOP LEVEL CELL: Or2Gate{sch}
XInverter@0 Out net@0 _16BitAdder__Inverter
XNor2Gate@0 net@0 Inp0 Inp1 _16BitAdder__Nor2Gate

* Spice Code nodes in cell cell 'Or2Gate{sch}'
vdd Vdd 0 DC 5
vin Inp0 0 DC 5 pulse(0 5 10f 0.5f 0.5f 20n 40n)
vin2 Inp1 0 DC 5 pulse(0 5 10f 0.5f 0.5f 40n 80n)
cload Out 0 50fF
.tran 0 100ns
.include C5_models.txt
.END
.END
