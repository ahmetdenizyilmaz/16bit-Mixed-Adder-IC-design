*** SPICE deck for cell 16BitMixedAdder{lay} from library 16BitAdder
*** Created on Sal Oca 08, 2019 18:54:37
*** Last revised on Paz Oca 13, 2019 23:12:13
*** Written on Pzt Oca 14, 2019 01:32:23 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT _16BitAdder__Inverter FROM CELL Inverter{lay}
.SUBCKT _16BitAdder__Inverter gnd Out vdd Inp
Mnmos@0 Out Inp gnd gnd NMOS L=0.6U W=1.8U AS=5.22P AD=4.455P PS=12.9U PD=8.7U
Mpmos@0 Out Inp vdd vdd PMOS L=0.6U W=3.6U AS=8.19P AD=4.455P PS=16.5U PD=8.7U
.ENDS _16BitAdder__Inverter

*** SUBCIRCUIT _16BitAdder__Nand2Gate FROM CELL Nand2Gate{lay}
.SUBCKT _16BitAdder__Nand2Gate gnd Out vdd Inp0 Inp1
Mnmos@0 net@32 Inp0 gnd gnd NMOS L=0.6U W=3.6U AS=8.19P AD=1.89P PS=16.5U PD=5.1U
Mnmos@1 Out Inp1 net@32 gnd NMOS L=0.6U W=3.6U AS=1.89P AD=4.14P PS=5.1U PD=7.1U
Mpmos@0 vdd Inp1 Out vdd PMOS L=0.6U W=3.6U AS=4.14P AD=7.065P PS=7.1U PD=13.5U
Mpmos@1 Out Inp0 vdd vdd PMOS L=0.6U W=3.6U AS=7.065P AD=4.14P PS=13.5U PD=7.1U
.ENDS _16BitAdder__Nand2Gate

*** SUBCIRCUIT _16BitAdder__And2Gate FROM CELL And2Gate{lay}
.SUBCKT _16BitAdder__And2Gate gnd Out vdd Inp0 Inp1
XInverter@0 gnd Out vdd net@2 _16BitAdder__Inverter
XNand2Gat@0 gnd net@2 vdd Inp0 Inp1 _16BitAdder__Nand2Gate
.ENDS _16BitAdder__And2Gate

*** SUBCIRCUIT _16BitAdder__Nor2Gate FROM CELL Nor2Gate{lay}
.SUBCKT _16BitAdder__Nor2Gate gnd Out vdd Inp0 Inp1
Mnmos@0 Out Inp0 gnd gnd NMOS L=0.6U W=1.8U AS=4.095P AD=3.06P PS=9.9U PD=5.9U
Mnmos@1 gnd Inp1 Out gnd NMOS L=0.6U W=1.8U AS=3.06P AD=4.095P PS=5.9U PD=9.9U
Mpmos@0 net@24 Inp0 vdd vdd PMOS L=0.6U W=3.6U AS=8.19P AD=2.025P PS=16.5U PD=5.4U
Mpmos@1 Out Inp1 net@24 vdd PMOS L=0.6U W=3.6U AS=2.025P AD=3.06P PS=5.4U PD=5.9U
.ENDS _16BitAdder__Nor2Gate

*** SUBCIRCUIT _16BitAdder__Or2Gate FROM CELL Or2Gate{lay}
.SUBCKT _16BitAdder__Or2Gate gnd Out vdd Inp0 Inp1
XInverter@2 gnd Out vdd net@8 _16BitAdder__Inverter
XNor2Gate@0 gnd net@8 vdd Inp0 Inp1 _16BitAdder__Nor2Gate
.ENDS _16BitAdder__Or2Gate

*** SUBCIRCUIT _16BitAdder__XorGate FROM CELL XorGate{lay}
.SUBCKT _16BitAdder__XorGate gnd Out vdd Inp0 Inp1
XNand2Gat@0 gnd net@17 vdd Inp0 Inp1 _16BitAdder__Nand2Gate
XNand2Gat@1 gnd net@23 vdd Inp0 net@17 _16BitAdder__Nand2Gate
XNand2Gat@4 gnd net@27 vdd net@17 Inp1 _16BitAdder__Nand2Gate
XNand2Gat@5 gnd Out vdd net@23 net@27 _16BitAdder__Nand2Gate
.ENDS _16BitAdder__XorGate

*** SUBCIRCUIT _16BitAdder__1BitAdder FROM CELL 1BitAdder{lay}
.SUBCKT _16BitAdder__1BitAdder Cin G0 gnd P0 Sum vdd Inp0 Inp1
XAnd2Gate@0 gnd G0 vdd Inp0 Inp1 _16BitAdder__And2Gate
XOr2Gate@0 gnd P0 vdd Inp0 Inp1 _16BitAdder__Or2Gate
XXorGate@0 gnd net@2 vdd Inp0 Inp1 _16BitAdder__XorGate
XXorGate@1 gnd Sum vdd net@2 Cin _16BitAdder__XorGate
.ENDS _16BitAdder__1BitAdder

*** SUBCIRCUIT _16BitAdder__CLAblock FROM CELL CLAblock{lay}
.SUBCKT _16BitAdder__CLAblock ChOut ClInp GhlOut GhInp GlInp gnd PhlOut PhInp PlInp vdd
XAnd2Gate@0 gnd PhlOut vdd PhInp PlInp _16BitAdder__And2Gate
XAnd2Gate@1 gnd net@39 vdd PhInp GlInp _16BitAdder__And2Gate
XAnd2Gate@2 gnd And2Gate@2_Out vdd ClInp PlInp _16BitAdder__And2Gate
XOr2Gate@1 gnd Or2Gate@1_Out vdd GhInp net@39 _16BitAdder__Or2Gate
XOr2Gate@2 gnd Or2Gate@2_Out vdd Or2Gate@2_Inp0 GlInp _16BitAdder__Or2Gate
.ENDS _16BitAdder__CLAblock

*** SUBCIRCUIT _16BitAdder__8BitCLAadder FROM CELL 8BitCLAadder{lay}
.SUBCKT _16BitAdder__8BitCLAadder A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 Cin gnd S0 S1 S2 S3 S4 S5 S6 S7 vdd
X_1BitAdde@0 net@5 net@0 gnd net@4 S7 vdd B7 A7 _16BitAdder__1BitAdder
X_1BitAdde@1 net@7 net@22 gnd net@15 S6 vdd B6 A6 _16BitAdder__1BitAdder
X_1BitAdde@2 net@50 net@52 gnd net@51 S5 vdd B5 A5 _16BitAdder__1BitAdder
X_1BitAdde@3 net@11 net@80 gnd net@87 S4 vdd B4 A4 _16BitAdder__1BitAdder
X_1BitAdde@4 net@527 net@128 gnd net@129 S3 vdd B3 A3 _16BitAdder__1BitAdder
X_1BitAdde@5 net@184 net@171 gnd net@176 S2 vdd B2 A2 _16BitAdder__1BitAdder
X_1BitAdde@6 net@225 net@221 gnd net@222 S1 vdd B1 A1 _16BitAdder__1BitAdder
X_1BitAdde@7 Cin net@250 gnd net@264 S0 vdd B0 A0 _16BitAdder__1BitAdder
XCLAblock@0 net@5 net@7 net@9 net@0 net@22 gnd net@8 net@4 net@15 vdd _16BitAdder__CLAblock
XCLAblock@1 net@7 net@11 net@12 net@9 net@66 gnd net@10 net@8 net@59 vdd _16BitAdder__CLAblock
XCLAblock@2 net@11 Cin CLAblock@2_GhlOut net@12 net@134 gnd CLAblock@2_PhlOut net@10 net@141 vdd _16BitAdder__CLAblock
XCLAblock@3 net@50 net@11 net@66 net@52 net@80 gnd net@59 net@51 net@87 vdd _16BitAdder__CLAblock
XCLAblock@4 net@527 net@184 net@131 net@128 net@171 gnd net@132 net@129 net@176 vdd _16BitAdder__CLAblock
XCLAblock@5 net@184 Cin net@134 net@131 net@227 gnd net@141 net@132 net@230 vdd _16BitAdder__CLAblock
XCLAblock@6 net@225 Cin net@227 net@221 net@250 gnd net@230 net@222 net@264 vdd _16BitAdder__CLAblock
.ENDS _16BitAdder__8BitCLAadder

*** SUBCIRCUIT _16BitAdder__Nand3Gate FROM CELL Nand3Gate{lay}
.SUBCKT _16BitAdder__Nand3Gate gnd Out vdd Inp0 Inp1 Inp2
Mnmos@0 Out Inp2 net@18 gnd NMOS L=0.6U W=5.4U AS=2.7P AD=5.333P PS=6.9U PD=8.85U
Mnmos@1 net@19 Inp0 gnd gnd NMOS L=0.6U W=5.4U AS=11.16P AD=2.835P PS=20.1U PD=7.2U
Mnmos@2 net@18 Inp1 net@19 gnd NMOS L=0.6U W=5.4U AS=2.835P AD=2.7P PS=7.2U PD=6.9U
Mpmos@0 Out Inp2 vdd vdd PMOS L=0.6U W=3.6U AS=5.04P AD=5.333P PS=9.3U PD=8.85U
Mpmos@1 vdd Inp1 Out vdd PMOS L=0.6U W=3.6U AS=5.333P AD=5.04P PS=8.85U PD=9.3U
Mpmos@2 Out Inp0 vdd vdd PMOS L=0.6U W=3.6U AS=5.04P AD=5.333P PS=9.3U PD=8.85U
.ENDS _16BitAdder__Nand3Gate

*** SUBCIRCUIT _16BitAdder__1BitFA FROM CELL 1BitFA{lay}
.SUBCKT _16BitAdder__1BitFA Cin Cout gnd Sum Testand1 Testand2 Testand3 vdd Inp0 Inp1
XNand2Gat@0 gnd Testand1 vdd Inp0 Inp1 _16BitAdder__Nand2Gate
XNand2Gat@1 gnd Testand2 vdd Cin Inp1 _16BitAdder__Nand2Gate
XNand2Gat@2 gnd Testand3 vdd Cin Inp0 _16BitAdder__Nand2Gate
XNand3Gat@0 gnd Cout vdd Testand1 Testand2 Testand3 _16BitAdder__Nand3Gate
XXorGate@0 gnd net@90 vdd Inp0 Inp1 _16BitAdder__XorGate
XXorGate@1 gnd Sum vdd net@90 Cin _16BitAdder__XorGate
.ENDS _16BitAdder__1BitFA

*** SUBCIRCUIT _16BitAdder__4bitFA FROM CELL 4bitFA{lay}
.SUBCKT _16BitAdder__4bitFA A0 A1 A2 A3 B0 B1 B2 B3 Cin Cout gnd S0 S1 S2 S3 vdd
X_1BitFA@0 net@2 net@0 gnd S2 _1BitFA@0_Testand1 _1BitFA@0_Testand2 _1BitFA@0_Testand3 vdd A2 B2 _16BitAdder__1BitFA
X_1BitFA@1 net@0 Cout gnd S3 _1BitFA@1_Testand1 _1BitFA@1_Testand2 _1BitFA@1_Testand3 vdd A3 B3 _16BitAdder__1BitFA
X_1BitFA@2 net@1 net@2 gnd S1 _1BitFA@2_Testand1 _1BitFA@2_Testand2 _1BitFA@2_Testand3 vdd A1 B1 _16BitAdder__1BitFA
X_1BitFA@3 Cin net@1 gnd S0 _1BitFA@3_Testand1 _1BitFA@3_Testand2 _1BitFA@3_Testand3 vdd A0 B0 _16BitAdder__1BitFA
.ENDS _16BitAdder__4bitFA

*** SUBCIRCUIT _16BitAdder__8BitFA FROM CELL 8BitFA{lay}
.SUBCKT _16BitAdder__8BitFA A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 Cin Cout GND S0 S1 S2 S3 S4 S5 S6 S7 vdd
X_4bitFA@0 A4 A5 A6 A7 B4 B5 B6 B7 net@0 Cout GND S4 S5 S6 S7 vdd _16BitAdder__4bitFA
X_4bitFA@1 A0 A1 A2 A3 B0 B1 B2 B3 Cin net@0 GND S0 S1 S2 S3 vdd _16BitAdder__4bitFA
.ENDS _16BitAdder__8BitFA

*** TOP LEVEL CELL: 16BitMixedAdder{lay}
X_8BitCLAa@0 A8 A9 A10 A11 A12 A13 A14 A15 B8 B9 B10 B11 B12 B13 B14 B15 net@0 gnd S8 S9 S10 S11 S12 S13 S14 S15 vdd _16BitAdder__8BitCLAadder
X_8BitFA@0 A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 Cin net@0 gnd S0 S1 S2 S3 S4 S5 S6 S7 vdd _16BitAdder__8BitFA

* Spice Code nodes in cell cell '16BitMixedAdder{lay}'

vdd Vdd 0 DC 5
vin A0 0 DC 0
vin2 A1 0 DC 5
vin3 A2 0 DC 5
vin4 A3 0 DC 5
vin5 A4 0 DC 5
vin6 A5 0 DC 5
vin7 A6 0 DC 5
vin8 A7 0 DC 5
vin9 A8 0 DC 0
vin10 A9 0 DC 0
vin11 A10 0 DC 0
vin12 A11 0 DC 0
vin13 A12 0 DC 0
vin14 A13 0 DC 0
vin15 A14 0 DC 0
vin16 A15 0 DC 0

vin17 B0 0 DC 0
vin18 B1 0 DC 0
vin19 B2 0 DC 0
vin20 B3 0 DC 0
vin21 B4 0 DC 0
vin22 B5 0 DC 0
vin23 B6 0 DC 0
vin24 B7 0 DC 0
vin25 B8 0 DC 0
vin26 B9 0 DC 0
vin27 B10 0 DC 0
vin28 B11 0 DC 0
vin29 B12 0 DC 0
vin30 B13 0 DC 0
vin31 B14 0 DC 5
vin32 B15 0 DC 0

.tran 10ns 100ns
.include C5_models.txt
.END
.END
