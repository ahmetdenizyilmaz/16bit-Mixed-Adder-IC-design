*** SPICE deck for cell And2Gate{sch} from library 16BitAdder
*** Created on Pzt Oca 07, 2019 17:56:27
*** Last revised on Paz Oca 13, 2019 20:31:54
*** Written on Paz Oca 13, 2019 20:31:56 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT _16BitAdder__Inverter FROM CELL Inverter{sch}
.SUBCKT _16BitAdder__Inverter Out Inp
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 Out Inp gnd gnd NMOS L=0.6U W=1.8U
Mpmos@1 vdd Inp Out vdd PMOS L=0.6U W=3.6U
.ENDS _16BitAdder__Inverter

*** SUBCIRCUIT _16BitAdder__Nand2Gate FROM CELL Nand2Gate{sch}
.SUBCKT _16BitAdder__Nand2Gate Out Inp0 Inp1
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@1 Inp1 gnd gnd NMOS L=0.6U W=3.6U
Mnmos@1 Out Inp0 net@1 gnd NMOS L=0.6U W=3.6U
Mpmos@0 vdd Inp1 Out vdd PMOS L=0.6U W=3.6U
Mpmos@1 vdd Inp0 Out vdd PMOS L=0.6U W=3.6U
.ENDS _16BitAdder__Nand2Gate

.global gnd vdd

*** TOP LEVEL CELL: And2Gate{sch}
XInverter@1 Out net@8 _16BitAdder__Inverter
XNand2Gat@0 net@8 Inp0 Inp1 _16BitAdder__Nand2Gate

* Spice Code nodes in cell cell 'And2Gate{sch}'
vdd Vdd 0 DC 5
vin Inp0 0 DC 5 pulse(0 5 10f 0.5f 0.5f 20n 40n)
vin2 Inp1 0 DC 5 pulse(0 5 10f 0.5f 0.5f 40n 80n)
cload Out 0 50fF
.tran 0 100ns
.include C5_models.txt
.END
.END
