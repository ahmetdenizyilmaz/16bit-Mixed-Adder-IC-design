*** SPICE deck for cell 8BitFA{sch} from library 16BitAdder
*** Created on Sal Oca 08, 2019 18:34:56
*** Last revised on Paz Oca 13, 2019 22:07:10
*** Written on Paz Oca 13, 2019 22:09:58 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT _16BitAdder__Nand2Gate FROM CELL Nand2Gate{sch}
.SUBCKT _16BitAdder__Nand2Gate Out Inp0 Inp1
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@1 Inp1 gnd gnd NMOS L=0.6U W=3.6U
Mnmos@1 Out Inp0 net@1 gnd NMOS L=0.6U W=3.6U
Mpmos@0 vdd Inp1 Out vdd PMOS L=0.6U W=3.6U
Mpmos@1 vdd Inp0 Out vdd PMOS L=0.6U W=3.6U
.ENDS _16BitAdder__Nand2Gate

*** SUBCIRCUIT _16BitAdder__Nand3Gate FROM CELL Nand3Gate{sch}
.SUBCKT _16BitAdder__Nand3Gate Out Inp0 Inp1 Inp2
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@20 Inp0 gnd gnd NMOS L=0.6U W=5.4U
Mnmos@1 net@21 Inp1 net@20 gnd NMOS L=0.6U W=5.4U
Mnmos@2 Out Inp2 net@21 gnd NMOS L=0.6U W=5.4U
Mpmos@0 vdd Inp0 Out vdd PMOS L=0.6U W=3.6U
Mpmos@1 vdd Inp1 Out vdd PMOS L=0.6U W=3.6U
Mpmos@2 vdd Inp2 Out vdd PMOS L=0.6U W=3.6U
.ENDS _16BitAdder__Nand3Gate

*** SUBCIRCUIT _16BitAdder__XorGate FROM CELL XorGate{sch}
.SUBCKT _16BitAdder__XorGate Out Inp0 Inp1
** GLOBAL gnd
** GLOBAL vdd
XNand2Gat@0 net@14 Inp0 net@0 _16BitAdder__Nand2Gate
XNand2Gat@1 net@15 net@0 Inp1 _16BitAdder__Nand2Gate
XNand2Gat@3 Out net@14 net@15 _16BitAdder__Nand2Gate
XNand2Gat@4 net@0 Inp0 Inp1 _16BitAdder__Nand2Gate
.ENDS _16BitAdder__XorGate

*** SUBCIRCUIT _16BitAdder__1BitFA FROM CELL 1BitFA{sch}
.SUBCKT _16BitAdder__1BitFA Cin Cout Sum Inp0 Inp1
** GLOBAL gnd
** GLOBAL vdd
XNand2Gat@0 net@0 Inp0 Inp1 _16BitAdder__Nand2Gate
XNand2Gat@1 net@2 Inp0 Cin _16BitAdder__Nand2Gate
XNand2Gat@2 net@3 Inp1 Cin _16BitAdder__Nand2Gate
XNand3Gat@0 Cout net@0 net@2 net@3 _16BitAdder__Nand3Gate
XXorGate@0 net@8 Inp0 Inp1 _16BitAdder__XorGate
XXorGate@1 Sum net@8 Cin _16BitAdder__XorGate
.ENDS _16BitAdder__1BitFA

*** SUBCIRCUIT _16BitAdder__4bitFA FROM CELL 4bitFA{sch}
.SUBCKT _16BitAdder__4bitFA A0 A1 A2 A3 B0 B1 B2 B3 Cin Cout S0 S1 S2 S3
** GLOBAL gnd
** GLOBAL vdd
Rres@2 gnd Cin 100k
X_1BitFA@8 net@52 Cout S3 A3 B3 _16BitAdder__1BitFA
X_1BitFA@9 net@57 net@52 S2 A2 B2 _16BitAdder__1BitFA
X_1BitFA@10 net@64 net@57 S1 A1 B1 _16BitAdder__1BitFA
X_1BitFA@11 Cin net@64 S0 A0 B0 _16BitAdder__1BitFA
.ENDS _16BitAdder__4bitFA

.global gnd vdd

*** TOP LEVEL CELL: 8BitFA{sch}
X_4bitFA@0 A0 A1 A2 A3 B0 B1 B2 B3 _4bitFA@0_Cin net@1 S0 S1 S2 S3 _16BitAdder__4bitFA
X_4bitFA@1 A4 A5 A6 A7 B4 B5 B6 B7 net@1 _4bitFA@1_Cout S4 S5 S6 S7 _16BitAdder__4bitFA

* Spice Code nodes in cell cell '8BitFA{sch}'
vdd Vdd 0 DC 5

vin A0 0 DC 5
vin2 A1 0 DC 0
vin3 A2 0 DC 5
vin4 A3 0 DC 0
vin5 A4 0 DC 5
vin6 A5 0 DC 5
vin7 A6 0 DC 0
vin8 A7 0 DC 0

vin9 B0 0 DC 5
vin10 B1 0 DC 5
vin11 B2 0 DC 5
vin12 B3 0 DC 5
vin13 B4 0 DC 5
vin14 B5 0 DC 5
vin15 B6 0 DC 0
vin16 B7 0 DC 5

cload S0 0 5fF
.tran 0 100ns
.include C5_models.txt
.END
