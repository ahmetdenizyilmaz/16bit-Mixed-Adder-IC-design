*** SPICE deck for cell Nand2Gate{lay} from library Fulladder2
*** Created on Çar Ara 20, 2000 23:56:15
*** Last revised on Paz Oca 13, 2019 18:05:26
*** Written on Paz Oca 13, 2019 18:05:28 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: Nand2Gate{lay}
Mnmos@0 net@32 Inp0 gnd gnd NMOS L=0.6U W=3.6U AS=8.19P AD=1.89P PS=16.5U PD=5.1U
Mnmos@1 Out Inp1 net@32 gnd NMOS L=0.6U W=3.6U AS=1.89P AD=4.14P PS=5.1U PD=7.1U
Mpmos@0 vdd Inp1 Out vdd PMOS L=0.6U W=3.6U AS=4.14P AD=7.065P PS=7.1U PD=13.5U
Mpmos@1 Out Inp0 vdd vdd PMOS L=0.6U W=3.6U AS=7.065P AD=4.14P PS=13.5U PD=7.1U

* Spice Code nodes in cell cell 'Nand2Gate{lay}'
vdd Vdd 0 DC 5
vin Inp0 0 DC 5 pulse(0 5 10f 0.5f 0.5f 20n 40n)
vin2 Inp1 0 DC 5 pulse(0 5 10f 0.5f 0.5f 40n 80n)
cload Out 0 50fF
.tran 0 100ns
.include C5_models.txt
.END

