*** SPICE deck for cell 8BitCLAadder{sch} from library 16BitAdder
*** Created on Pzt Oca 07, 2019 20:17:35
*** Last revised on Paz Oca 13, 2019 22:47:37
*** Written on Paz Oca 13, 2019 22:57:21 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT _16BitAdder__Inverter FROM CELL Inverter{sch}
.SUBCKT _16BitAdder__Inverter Out Inp
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 Out Inp gnd gnd NMOS L=0.6U W=1.8U
Mpmos@1 vdd Inp Out vdd PMOS L=0.6U W=3.6U
.ENDS _16BitAdder__Inverter

*** SUBCIRCUIT _16BitAdder__Nand2Gate FROM CELL Nand2Gate{sch}
.SUBCKT _16BitAdder__Nand2Gate Out Inp0 Inp1
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@1 Inp1 gnd gnd NMOS L=0.6U W=3.6U
Mnmos@1 Out Inp0 net@1 gnd NMOS L=0.6U W=3.6U
Mpmos@0 vdd Inp1 Out vdd PMOS L=0.6U W=3.6U
Mpmos@1 vdd Inp0 Out vdd PMOS L=0.6U W=3.6U
.ENDS _16BitAdder__Nand2Gate

*** SUBCIRCUIT _16BitAdder__And2Gate FROM CELL And2Gate{sch}
.SUBCKT _16BitAdder__And2Gate Out Inp0 Inp1
** GLOBAL gnd
** GLOBAL vdd
XInverter@1 Out net@8 _16BitAdder__Inverter
XNand2Gat@0 net@8 Inp0 Inp1 _16BitAdder__Nand2Gate
.ENDS _16BitAdder__And2Gate

*** SUBCIRCUIT _16BitAdder__Nor2Gate FROM CELL Nor2Gate{sch}
.SUBCKT _16BitAdder__Nor2Gate Out Inp0 Inp1
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Out Inp0 gnd gnd NMOS L=0.6U W=1.8U
Mnmos@1 Out Inp1 gnd gnd NMOS L=0.6U W=1.8U
Mpmos@0 net@11 Inp1 Out vdd PMOS L=0.6U W=3.6U
Mpmos@1 vdd Inp0 net@11 vdd PMOS L=0.6U W=3.6U
.ENDS _16BitAdder__Nor2Gate

*** SUBCIRCUIT _16BitAdder__Or2Gate FROM CELL Or2Gate{sch}
.SUBCKT _16BitAdder__Or2Gate Out Inp0 Inp1
** GLOBAL gnd
** GLOBAL vdd
XInverter@0 Out net@0 _16BitAdder__Inverter
XNor2Gate@0 net@0 Inp0 Inp1 _16BitAdder__Nor2Gate
.ENDS _16BitAdder__Or2Gate

*** SUBCIRCUIT _16BitAdder__XorGate FROM CELL XorGate{sch}
.SUBCKT _16BitAdder__XorGate Out Inp0 Inp1
** GLOBAL gnd
** GLOBAL vdd
XNand2Gat@0 net@14 Inp0 net@0 _16BitAdder__Nand2Gate
XNand2Gat@1 net@15 net@0 Inp1 _16BitAdder__Nand2Gate
XNand2Gat@3 Out net@14 net@15 _16BitAdder__Nand2Gate
XNand2Gat@4 net@0 Inp0 Inp1 _16BitAdder__Nand2Gate
.ENDS _16BitAdder__XorGate

*** SUBCIRCUIT _16BitAdder__1BitAdder FROM CELL 1BitAdder{sch}
.SUBCKT _16BitAdder__1BitAdder Cin G0 P0 Sum Inp0 Inp1
** GLOBAL gnd
** GLOBAL vdd
XAnd2Gate@0 G0 Inp0 Inp1 _16BitAdder__And2Gate
XOr2Gate@0 P0 Inp0 Inp1 _16BitAdder__Or2Gate
XXorGate@0 net@13 Inp0 Inp1 _16BitAdder__XorGate
XXorGate@1 Sum net@13 Cin _16BitAdder__XorGate
.ENDS _16BitAdder__1BitAdder

*** SUBCIRCUIT _16BitAdder__CLAblock FROM CELL CLAblock{sch}
.SUBCKT _16BitAdder__CLAblock ChOut ClInp GhlOut GhInp GlInp PhlOut PhInp PlInp
** GLOBAL gnd
** GLOBAL vdd
XAnd2Gate@0 PhlOut PlInp PhInp _16BitAdder__And2Gate
XAnd2Gate@1 net@4 GlInp And2Gate@1_Inp1 _16BitAdder__And2Gate
XAnd2Gate@2 net@18 ClInp PlInp _16BitAdder__And2Gate
XOr2Gate@0 GhlOut net@4 GhInp _16BitAdder__Or2Gate
XOr2Gate@1 ChOut net@18 GlInp _16BitAdder__Or2Gate
.ENDS _16BitAdder__CLAblock

.global gnd vdd

*** TOP LEVEL CELL: 8BitCLAadder{sch}
X_1BitAdde@0 net@2 net@0 net@1 S7 A7 B7 _16BitAdder__1BitAdder
X_1BitAdde@1 net@5 net@9 net@11 S6 A6 B6 _16BitAdder__1BitAdder
X_1BitAdde@2 net@17 net@15 net@16 S5 A5 B5 _16BitAdder__1BitAdder
X_1BitAdde@3 net@8 net@24 net@26 S4 A4 B4 _16BitAdder__1BitAdder
X_1BitAdde@4 net@32 net@30 net@31 S3 A3 B3 _16BitAdder__1BitAdder
X_1BitAdde@5 net@37 net@33 net@35 S2 A2 B2 _16BitAdder__1BitAdder
X_1BitAdde@6 net@45 net@43 net@44 S1 A1 B1 _16BitAdder__1BitAdder
X_1BitAdde@7 Cin net@52 net@54 S0 A0 B0 _16BitAdder__1BitAdder
XCLAblock@0 net@2 net@5 net@3 net@0 net@9 net@4 net@1 net@11 _16BitAdder__CLAblock
XCLAblock@1 net@5 net@8 net@6 net@3 net@18 net@7 net@4 net@20 _16BitAdder__CLAblock
XCLAblock@2 net@8 Cin CLAblock@2_GhlOut net@6 net@58 CLAblock@2_PhlOut net@7 net@60 _16BitAdder__CLAblock
XCLAblock@3 net@17 net@8 net@18 net@15 net@24 net@20 net@16 net@26 _16BitAdder__CLAblock
XCLAblock@4 net@32 net@37 net@40 net@30 net@33 net@41 net@31 net@35 _16BitAdder__CLAblock
XCLAblock@5 net@37 Cin net@58 net@40 net@46 net@60 net@41 net@48 _16BitAdder__CLAblock
XCLAblock@6 net@45 Cin net@46 net@43 net@52 net@48 net@44 net@54 _16BitAdder__CLAblock

* Spice Code nodes in cell cell '8BitCLAadder{sch}'
vvdd Vdd 0 DC 5
*A Bits
vin A0 0 DC 5
vin2 A1 0 DC 5
vin3 A2 0 DC 0
vin4 A3 0 DC 5
vin5 A4 0 DC 5
vin6 A5 0 DC 0
vin7 A6 0 DC 5
vin8 A7 0 DC 5
*B Bits
vin9 B0 0 DC 0
vin10 B1 0 DC 5
vin11 B2 0 DC 0
vin12 B3 0 DC 0
vin13 B4 0 DC 5
vin14 B5 0 DC 0
vin15 B6 0 DC 0
vin16 B7 0 DC 0
cload S0 0 5fF
.tran 0 100ns
.include C5_models.txt
.END

