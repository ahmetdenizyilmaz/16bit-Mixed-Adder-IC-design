*** SPICE deck for cell 1BitFA{lay} from library 16BitAdder
*** Created on Pzt Oca 07, 2019 00:37:02
*** Last revised on Paz Oca 13, 2019 21:35:40
*** Written on Paz Oca 13, 2019 21:35:46 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT _16BitAdder__Nand2Gate FROM CELL Nand2Gate{lay}
.SUBCKT _16BitAdder__Nand2Gate gnd Out vdd Inp0 Inp1
Mnmos@0 net@32 Inp0 gnd gnd NMOS L=0.6U W=3.6U AS=8.19P AD=1.89P PS=16.5U PD=5.1U
Mnmos@1 Out Inp1 net@32 gnd NMOS L=0.6U W=3.6U AS=1.89P AD=4.14P PS=5.1U PD=7.1U
Mpmos@0 vdd Inp1 Out vdd PMOS L=0.6U W=3.6U AS=4.14P AD=7.065P PS=7.1U PD=13.5U
Mpmos@1 Out Inp0 vdd vdd PMOS L=0.6U W=3.6U AS=7.065P AD=4.14P PS=13.5U PD=7.1U
.ENDS _16BitAdder__Nand2Gate

*** SUBCIRCUIT _16BitAdder__Nand3Gate FROM CELL Nand3Gate{lay}
.SUBCKT _16BitAdder__Nand3Gate gnd Out vdd Inp0 Inp1 Inp2
Mnmos@0 Out Inp2 net@18 gnd NMOS L=0.6U W=5.4U AS=2.7P AD=5.333P PS=6.9U PD=8.85U
Mnmos@1 net@19 Inp0 gnd gnd NMOS L=0.6U W=5.4U AS=11.16P AD=2.835P PS=20.1U PD=7.2U
Mnmos@2 net@18 Inp1 net@19 gnd NMOS L=0.6U W=5.4U AS=2.835P AD=2.7P PS=7.2U PD=6.9U
Mpmos@0 Out Inp2 vdd vdd PMOS L=0.6U W=3.6U AS=5.04P AD=5.333P PS=9.3U PD=8.85U
Mpmos@1 vdd Inp1 Out vdd PMOS L=0.6U W=3.6U AS=5.333P AD=5.04P PS=8.85U PD=9.3U
Mpmos@2 Out Inp0 vdd vdd PMOS L=0.6U W=3.6U AS=5.04P AD=5.333P PS=9.3U PD=8.85U
.ENDS _16BitAdder__Nand3Gate

*** SUBCIRCUIT _16BitAdder__XorGate FROM CELL XorGate{lay}
.SUBCKT _16BitAdder__XorGate gnd Out vdd Inp0 Inp1
XNand2Gat@0 gnd net@17 vdd Inp0 Inp1 _16BitAdder__Nand2Gate
XNand2Gat@1 gnd net@23 vdd Inp0 net@17 _16BitAdder__Nand2Gate
XNand2Gat@4 gnd net@27 vdd net@17 Inp1 _16BitAdder__Nand2Gate
XNand2Gat@5 gnd Out vdd net@23 net@27 _16BitAdder__Nand2Gate
.ENDS _16BitAdder__XorGate

*** TOP LEVEL CELL: 1BitFA{lay}
XNand2Gat@0 gnd Testand1 vdd Inp0 Inp1 _16BitAdder__Nand2Gate
XNand2Gat@1 gnd Testand2 vdd Cin Inp1 _16BitAdder__Nand2Gate
XNand2Gat@2 gnd Testand3 vdd Cin Inp0 _16BitAdder__Nand2Gate
XNand3Gat@0 gnd Cout vdd Testand1 Testand2 Testand3 _16BitAdder__Nand3Gate
XXorGate@0 gnd net@90 vdd Inp0 Inp1 _16BitAdder__XorGate
XXorGate@1 gnd Sum vdd net@90 Cin _16BitAdder__XorGate

* Spice Code nodes in cell cell '1BitFA{lay}'
vdd Vdd 0 DC 5
vin Inp0 0 DC 5 pulse(0 5 10f 0.5f 0.5f 10n 20n)
vin2 Inp1 0 DC 5 pulse(0 5 10f 0.5f 0.5f 20n 40n)
vin3 Cin 0 DC pulse(5 0 10f 0.5f 0.5f 40n 80n)
cload Sum 0 50fF
.tran 100ns
.include C5_models.txt
.END
