*** SPICE deck for cell 1BitFA{sch} from library 16BitAdder
*** Created on Pzt Oca 07, 2019 00:25:43
*** Last revised on Paz Oca 13, 2019 21:07:55
*** Written on Paz Oca 13, 2019 21:23:08 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT _16BitAdder__Nand2Gate FROM CELL Nand2Gate{sch}
.SUBCKT _16BitAdder__Nand2Gate Out Inp0 Inp1
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@1 Inp1 gnd gnd NMOS L=0.6U W=3.6U
Mnmos@1 Out Inp0 net@1 gnd NMOS L=0.6U W=3.6U
Mpmos@0 vdd Inp1 Out vdd PMOS L=0.6U W=3.6U
Mpmos@1 vdd Inp0 Out vdd PMOS L=0.6U W=3.6U
.ENDS _16BitAdder__Nand2Gate

*** SUBCIRCUIT _16BitAdder__Nand3Gate FROM CELL Nand3Gate{sch}
.SUBCKT _16BitAdder__Nand3Gate Out Inp0 Inp1 Inp2
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@20 Inp0 gnd gnd NMOS L=0.6U W=5.4U
Mnmos@1 net@21 Inp1 net@20 gnd NMOS L=0.6U W=5.4U
Mnmos@2 Out Inp2 net@21 gnd NMOS L=0.6U W=5.4U
Mpmos@0 vdd Inp0 Out vdd PMOS L=0.6U W=3.6U
Mpmos@1 vdd Inp1 Out vdd PMOS L=0.6U W=3.6U
Mpmos@2 vdd Inp2 Out vdd PMOS L=0.6U W=3.6U
.ENDS _16BitAdder__Nand3Gate

*** SUBCIRCUIT _16BitAdder__XorGate FROM CELL XorGate{sch}
.SUBCKT _16BitAdder__XorGate Out Inp0 Inp1
** GLOBAL gnd
** GLOBAL vdd
XNand2Gat@0 net@14 Inp0 net@0 _16BitAdder__Nand2Gate
XNand2Gat@1 net@15 net@0 Inp1 _16BitAdder__Nand2Gate
XNand2Gat@3 Out net@14 net@15 _16BitAdder__Nand2Gate
XNand2Gat@4 net@0 Inp0 Inp1 _16BitAdder__Nand2Gate
.ENDS _16BitAdder__XorGate

.global gnd vdd

*** TOP LEVEL CELL: 1BitFA{sch}
XNand2Gat@0 net@0 Inp0 Inp1 _16BitAdder__Nand2Gate
XNand2Gat@1 net@2 Inp0 Cin _16BitAdder__Nand2Gate
XNand2Gat@2 net@3 Inp1 Cin _16BitAdder__Nand2Gate
XNand3Gat@0 Cout net@0 net@2 net@3 _16BitAdder__Nand3Gate
XXorGate@0 net@8 Inp0 Inp1 _16BitAdder__XorGate
XXorGate@1 Sum net@8 Cin _16BitAdder__XorGate

* Spice Code nodes in cell cell '1BitFA{sch}'
vdd Vdd 0 DC 5
vin Inp0 0 DC 5 pulse(0 5 10f 0.5f 0.5f 10n 20n)
vin2 Inp1 0 DC 5 pulse(0 5 10f 0.5f 0.5f 20n 40n)
vin3 Cin 0 DC pulse(5 0 10f 0.5f 0.5f 40n 80n)
cload Sum 0 50fF
.tran 100ns
.include C5_models.txt
.END
.END
