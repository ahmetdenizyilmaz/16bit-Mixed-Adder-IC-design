*** SPICE deck for cell Nor2Gate{sch} from library 16BitAdder
*** Created on Pzt Oca 07, 2019 17:23:00
*** Last revised on Paz Oca 13, 2019 20:11:18
*** Written on Paz Oca 13, 2019 20:13:55 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: Nor2Gate{sch}
Mnmos@0 Out Inp0 gnd gnd NMOS L=0.6U W=1.8U
Mnmos@1 Out Inp1 gnd gnd NMOS L=0.6U W=1.8U
Mpmos@0 net@11 Inp1 Out vdd PMOS L=0.6U W=3.6U
Mpmos@1 vdd Inp0 net@11 vdd PMOS L=0.6U W=3.6U

* Spice Code nodes in cell cell 'Nor2Gate{sch}'
vdd Vdd 0 DC 5
vin Inp0 0 DC 5 pulse(0 5 10f 0.5f 0.5f 20n 40n)
vin2 Inp1 0 DC 5 pulse(0 5 10f 0.5f 0.5f 40n 80n)
cload Out 0 50fF
.tran 0 100ns
.include C5_models.txt
.END
.END
