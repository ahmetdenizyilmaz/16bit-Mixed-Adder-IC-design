*** SPICE deck for cell And2Gate{lay} from library 16BitAdder
*** Created on Pzt Oca 07, 2019 17:59:35
*** Last revised on Paz Oca 13, 2019 20:31:03
*** Written on Paz Oca 13, 2019 20:31:07 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT _16BitAdder__Inverter FROM CELL Inverter{lay}
.SUBCKT _16BitAdder__Inverter gnd Out vdd Inp
Mnmos@0 Out Inp gnd gnd NMOS L=0.6U W=1.8U AS=5.22P AD=4.455P PS=12.9U PD=8.7U
Mpmos@0 Out Inp vdd vdd PMOS L=0.6U W=3.6U AS=8.19P AD=4.455P PS=16.5U PD=8.7U
.ENDS _16BitAdder__Inverter

*** SUBCIRCUIT _16BitAdder__Nand2Gate FROM CELL Nand2Gate{lay}
.SUBCKT _16BitAdder__Nand2Gate gnd Out vdd Inp0 Inp1
Mnmos@0 net@32 Inp0 gnd gnd NMOS L=0.6U W=3.6U AS=8.19P AD=1.89P PS=16.5U PD=5.1U
Mnmos@1 Out Inp1 net@32 gnd NMOS L=0.6U W=3.6U AS=1.89P AD=4.14P PS=5.1U PD=7.1U
Mpmos@0 vdd Inp1 Out vdd PMOS L=0.6U W=3.6U AS=4.14P AD=7.065P PS=7.1U PD=13.5U
Mpmos@1 Out Inp0 vdd vdd PMOS L=0.6U W=3.6U AS=7.065P AD=4.14P PS=13.5U PD=7.1U
.ENDS _16BitAdder__Nand2Gate

*** TOP LEVEL CELL: And2Gate{lay}
XInverter@0 gnd Out vdd net@2 _16BitAdder__Inverter
XNand2Gat@0 gnd net@2 vdd Inp0 Inp1 _16BitAdder__Nand2Gate

* Spice Code nodes in cell cell 'And2Gate{lay}'
vdd Vdd 0 DC 5
vin Inp0 0 DC 5 pulse(0 5 10f 0.5f 0.5f 20n 40n)
vin2 Inp1 0 DC 5 pulse(0 5 10f 0.5f 0.5f 40n 80n)
cload Out 0 50fF
.tran 0 100ns
.include C5_models.txt
.END
.END
