*** SPICE deck for cell Or2Gate{lay} from library 16BitAdder
*** Created on Pzt Oca 07, 2019 17:34:04
*** Last revised on Paz Oca 13, 2019 20:54:54
*** Written on Paz Oca 13, 2019 20:54:57 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT _16BitAdder__Inverter FROM CELL Inverter{lay}
.SUBCKT _16BitAdder__Inverter gnd Out vdd Inp
Mnmos@0 Out Inp gnd gnd NMOS L=0.6U W=1.8U AS=5.22P AD=4.455P PS=12.9U PD=8.7U
Mpmos@0 Out Inp vdd vdd PMOS L=0.6U W=3.6U AS=8.19P AD=4.455P PS=16.5U PD=8.7U
.ENDS _16BitAdder__Inverter

*** SUBCIRCUIT _16BitAdder__Nor2Gate FROM CELL Nor2Gate{lay}
.SUBCKT _16BitAdder__Nor2Gate gnd Out vdd Inp0 Inp1
Mnmos@0 Out Inp0 gnd gnd NMOS L=0.6U W=1.8U AS=4.095P AD=3.06P PS=9.9U PD=5.9U
Mnmos@1 gnd Inp1 Out gnd NMOS L=0.6U W=1.8U AS=3.06P AD=4.095P PS=5.9U PD=9.9U
Mpmos@0 net@24 Inp0 vdd vdd PMOS L=0.6U W=3.6U AS=8.19P AD=2.025P PS=16.5U PD=5.4U
Mpmos@1 Out Inp1 net@24 vdd PMOS L=0.6U W=3.6U AS=2.025P AD=3.06P PS=5.4U PD=5.9U
.ENDS _16BitAdder__Nor2Gate

*** TOP LEVEL CELL: Or2Gate{lay}
XInverter@2 gnd Out vdd net@8 _16BitAdder__Inverter
XNor2Gate@0 gnd net@8 vdd Inp0 Inp1 _16BitAdder__Nor2Gate

* Spice Code nodes in cell cell 'Or2Gate{lay}'
vdd Vdd 0 DC 5
vin Inp0 0 DC 5 pulse(0 5 10f 0.5f 0.5f 20n 40n)
vin2 Inp1 0 DC 5 pulse(0 5 10f 0.5f 0.5f 40n 80n)
cload Out 0 50fF
.tran 100ns
.include C5_models.txt
.END
.END
